package f_parameters;	 
	parameter k = 13;
	parameter l = 6;
	parameter m1 = 16;
	parameter m2 = 1;
	parameter delay = k+l;
endpackage 