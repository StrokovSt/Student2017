package parameters;
parameter in = 8;
parameter regout = 16;
endpackage
